** sch_path: /home/nguyen2604/projects/CMOS_INVERTER/CMOS_INVERTER.sch
**.subckt CMOS_INVERTER
V1 vin GND PULSE(0 1.8 1ns 1ns 1ns 5ns 10ns)
vdd vdd GND 1.8
XM1 vout vin GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM2 vout vin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran 0.1n 100n
.save all
.control
	run
	plot v(Vin) v(Vout)
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.end
