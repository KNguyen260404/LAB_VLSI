magic
tech sky130A
timestamp 1762022522
<< nwell >>
rect 810 350 1100 515
<< nmos >>
rect 900 220 915 305
rect 1000 275 1015 305
rect 900 170 915 200
rect 1000 170 1015 250
<< pmos >>
rect 900 370 915 495
rect 1000 370 1015 495
<< ndiff >>
rect 850 300 900 305
rect 850 280 870 300
rect 890 280 900 300
rect 850 275 900 280
rect 850 220 900 250
rect 915 300 1000 305
rect 915 280 920 300
rect 940 280 970 300
rect 990 280 1000 300
rect 915 275 1000 280
rect 1015 300 1065 305
rect 1015 280 1020 300
rect 1040 280 1065 300
rect 1015 275 1065 280
rect 915 220 1000 250
rect 850 195 900 200
rect 850 175 870 195
rect 890 175 900 195
rect 850 170 900 175
rect 915 195 1000 200
rect 915 175 920 195
rect 940 175 970 195
rect 990 175 1000 195
rect 915 170 1000 175
rect 1015 220 1065 250
rect 1015 195 1065 200
rect 1015 175 1020 195
rect 1040 175 1065 195
rect 1015 170 1065 175
<< pdiff >>
rect 850 445 900 495
rect 850 440 870 445
rect 890 440 900 445
rect 850 415 900 420
rect 850 375 870 415
rect 890 375 900 415
rect 850 370 900 375
rect 915 445 1000 495
rect 915 440 920 445
rect 940 440 970 445
rect 990 440 1000 445
rect 915 415 1000 420
rect 915 375 920 415
rect 940 375 970 415
rect 990 375 1000 415
rect 915 370 1000 375
rect 1015 445 1065 495
rect 1015 440 1020 445
rect 1040 440 1065 445
rect 1015 415 1065 420
rect 1015 375 1020 415
rect 1040 375 1065 415
rect 1015 370 1065 375
<< ndiffc >>
rect 870 280 890 300
rect 920 280 940 300
rect 970 280 990 300
rect 1020 280 1040 300
rect 870 175 890 195
rect 920 175 940 195
rect 970 175 990 195
rect 1020 175 1040 195
<< pdiffc >>
rect 870 440 890 445
rect 870 375 890 415
rect 920 440 940 445
rect 970 440 990 445
rect 920 375 940 415
rect 970 375 990 415
rect 1020 440 1040 445
rect 1020 375 1040 415
<< psubdiff >>
rect 830 275 850 305
rect 830 220 850 250
rect 830 170 850 200
<< psubdiffcont >>
rect 830 250 850 275
<< nsubdiffcont >>
rect 830 375 850 415
<< poly >>
rect 900 495 915 510
rect 1000 495 1015 510
rect 900 305 915 370
rect 1000 305 1015 370
rect 1000 250 1015 275
rect 900 200 915 220
rect 900 155 915 170
rect 1000 155 1015 170
rect 875 150 915 155
rect 875 130 885 150
rect 905 130 915 150
rect 875 125 915 130
rect 975 150 1015 155
rect 975 130 985 150
rect 1005 130 1015 150
rect 975 125 1015 130
<< polycont >>
rect 815 520 825 530
rect 1000 520 1010 530
rect 885 130 905 150
rect 985 130 1005 150
<< locali >>
rect 850 440 870 445
rect 890 440 920 445
rect 940 440 970 445
rect 990 440 1020 445
rect 1040 440 1065 445
rect 1000 425 1010 440
rect 850 375 870 415
rect 890 375 920 415
rect 940 375 970 415
rect 990 375 1020 415
rect 1040 375 1065 415
rect 850 280 870 300
rect 890 280 920 300
rect 940 280 970 300
rect 990 280 1020 300
rect 1040 280 1065 300
rect 850 175 870 195
rect 890 175 920 195
rect 940 175 970 195
rect 990 175 1020 195
rect 1040 175 1065 195
rect 875 130 885 150
rect 975 130 985 150
<< viali >>
rect 815 450 825 520
rect 1000 445 1010 520
rect 870 440 890 445
rect 920 440 940 445
rect 970 440 990 445
rect 1020 440 1040 445
rect 870 425 890 440
rect 920 425 940 440
rect 970 425 990 440
rect 1020 425 1040 440
rect 830 375 850 415
rect 870 375 890 415
rect 920 375 940 415
rect 970 375 990 415
rect 1020 375 1040 415
rect 870 280 890 300
rect 920 280 940 300
rect 970 280 990 300
rect 1020 280 1040 300
rect 870 175 890 195
rect 920 175 940 195
rect 970 175 990 195
rect 1020 175 1040 195
<< metal1 >>
rect 810 450 815 490
rect 825 450 1000 490
rect 1010 450 1100 490
rect 810 425 870 445
rect 890 425 920 445
rect 940 425 970 445
rect 990 425 1020 445
rect 1040 425 1100 445
rect 810 375 830 415
rect 850 375 870 415
rect 890 375 920 415
rect 940 375 970 415
rect 990 375 1020 415
rect 1040 375 1100 415
rect 810 280 870 300
rect 890 280 920 300
rect 940 280 970 300
rect 990 280 1020 300
rect 1040 280 1100 300
rect 810 175 870 195
rect 890 175 920 195
rect 940 175 970 195
rect 990 175 1020 195
rect 1040 175 1100 195
rect 875 130 905 150
rect 975 130 1005 150
<< labels >>
rlabel metal1 810 140 810 140 7 A
port 1 w
rlabel metal1 1100 140 1100 140 3 B
port 2 e
rlabel metal1 1100 395 1100 395 3 Y
port 3 e
rlabel metal1 810 470 810 470 7 VDD
port 4 w
rlabel metal1 810 185 810 185 7 GND
port 5 w
<< end >>
