* SPICE3 file created from CMOS_NAND_test.ext - technology: sky130A

X0 VDD a_1750_250# Y Y sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.1 as=0.25 ps=2 w=1.05 l=0.15
X1 a_1700_550# a_1750_250# a_1700_440# a_1660_340# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.45 l=0.15
X2 VDD a_1950_250# Y Y sky130_fd_pr__pfet_01v8 ad=0.23375 pd=1.4 as=0.2125 ps=1.35 w=1.05 l=0.15
X3 GND a_1750_250# GND a_1660_340# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.555 ps=5.5 w=0.3 l=0.15
X4 a_1830_440# a_1950_250# GND a_1660_340# sky130_fd_pr__nfet_01v8 ad=0.1275 pd=1.15 as=0.1275 ps=1.15 w=0.45 l=0.15
X5 a_1700_550# a_1950_250# a_1700_550# a_1660_340# sky130_fd_pr__nfet_01v8 ad=0.1275 pd=1.15 as=0.555 ps=5.5 w=0.3 l=0.15
