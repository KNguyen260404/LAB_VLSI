** sch_path: /home/nguyen2604/projects/CMOS_NAND/CMOS_NAND_SCHEMATIC.sch
**.subckt CMOS_NAND_SCHEMATIC
XM1 Y A net1 net1 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM2 Y B VDD Y sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1 m=1
XM3 Y A VDD Y sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 B GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
V1 A GND PULSE(0 1.8 1.5n 10p 10p 50n 100n)
V2 VDD GND 1.8
V3 B GND PULSE(0 1.8 25n 10p 10p 50p 100n)
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran 0.1n 200n
.save all
.control
  run
  plot V(A) V(B) V(Y)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
