* SPICE3 file created from NMOS_TECH-ICC.ext - technology: sky130A

X0 a_1910_310# a_1880_280# a_1640_310# a_1640_310# sky130_fd_pr__nfet_01v8 ad=0.72 pd=3.6 as=0.72 ps=3.6 w=1.2 l=0.15
