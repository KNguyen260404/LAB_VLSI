magic
tech sky130A
timestamp 1762272601
<< error_p >>
rect 820 155 880 275
<< nmos >>
rect 940 155 955 275
<< ndiff >>
rect 880 255 940 275
rect 880 175 900 255
rect 920 175 940 255
rect 880 155 940 175
rect 955 255 1015 275
rect 955 175 975 255
rect 995 175 1015 255
rect 955 155 1015 175
<< ndiffc >>
rect 900 175 920 255
rect 975 175 995 255
<< psubdiff >>
rect 820 255 880 275
rect 820 175 840 255
rect 860 175 880 255
rect 820 155 880 175
<< psubdiffcont >>
rect 840 175 860 255
<< poly >>
rect 940 275 955 290
rect 940 140 955 155
<< locali >>
rect 825 255 935 270
rect 825 175 840 255
rect 860 175 900 255
rect 920 175 935 255
rect 825 160 935 175
rect 960 255 1010 270
rect 960 175 975 255
rect 995 175 1010 255
rect 960 160 1010 175
<< end >>
