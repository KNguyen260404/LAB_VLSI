** sch_path: /home/nguyen2604/projects/NMOS/NMOS.sch
**.subckt NMOS
XM1 net1 net2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
V1 net2 GND 0
V2 net1 GND 0.9
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.control
  dc V1 0 3 0.01
  plot -i(V2)
.endc
.save all


**** end user architecture code
**.ends
.GLOBAL GND
.end
