magic
tech sky130A
timestamp 1762022523
<< nwell >>
rect 810 350 1100 515
<< pmos >>
rect 900 420 915 440
rect 1000 420 1015 440
<< nmos >>
rect 900 250 915 275
rect 1000 200 1015 220
<< pdiff >>
rect 850 440 1065 495
rect 850 370 1065 420
<< ndiff >>
rect 850 275 1065 305
rect 850 220 1065 250
rect 850 170 1065 200
<< pdiffc >>
rect 870 450 890 490
rect 920 450 940 490
rect 970 450 990 490
rect 1020 450 1040 490
rect 870 375 890 415
rect 920 375 940 415
rect 970 375 990 415
rect 1020 375 1040 415
<< ndiffc >>
rect 870 280 890 300
rect 920 280 940 300
rect 970 280 990 300
rect 1020 280 1040 300
rect 870 175 890 195
rect 920 175 940 195
rect 970 175 990 195
rect 1020 175 1040 195
<< psubdiff >>
rect 830 275 850 305
rect 830 220 850 250
rect 830 170 850 200
<< nsubdiff >>
rect 830 440 850 495
rect 830 370 850 420
<< psubdiffcont >>
rect 830 250 850 275
<< nsubdiffcont >>
rect 830 440 850 495
<< poly >>
rect 900 155 915 510
rect 1000 155 1015 510
rect 875 125 915 155
rect 975 125 1015 155
<< polycont >>
rect 885 130 905 150
rect 985 130 1005 150
<< locali >>
rect 850 450 1065 490
rect 850 375 1065 415
rect 850 280 1065 300
rect 850 175 1065 195
rect 875 130 905 150
rect 975 130 1005 150
<< viali >>
rect 870 450 890 490
rect 920 450 940 490
rect 970 450 990 490
rect 1020 450 1040 490
rect 870 375 890 415
rect 920 375 940 415
rect 970 375 990 415
rect 1020 375 1040 415
rect 870 280 890 300
rect 920 280 940 300
rect 970 280 990 300
rect 1020 280 1040 300
rect 870 175 890 195
rect 920 175 940 195
rect 970 175 990 195
rect 1020 175 1040 195
<< metal1 >>
rect 810 450 1100 490
rect 810 375 1100 415
rect 810 280 1100 300
rect 810 175 1100 195
rect 875 130 905 150
rect 975 130 1005 150
<< labels >>
rlabel metal1 810 140 810 140 7 A
port 1 w
rlabel metal1 1100 140 1100 140 3 B
port 2 e
rlabel metal1 1100 395 1100 395 3 Y
port 3 e
rlabel metal1 810 470 810 470 7 VDD
port 4 w
rlabel metal1 810 185 810 185 7 GND
port 5 w
<< end >>

