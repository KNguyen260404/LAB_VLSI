M1 N006 N003 N005 0 myNMOS l=1u w=20u
M2 Vout N002 N005 0 myNMOS l=1u w=20u
M3 N004 N004 0 0 myNMOS l=1u w=10u
M4 N005 N004 0 0 myNMOS l=1u w=10u
M5 N001 N007 N006 N001 myPMOS l=0.5u w=20u
M6 N001 N007 N007 N001 myPMOS l=0.5u w=20u
M7 N001 N007 Vout N001 myPMOS l=0.5u w=20u
M8 Vout N004 0 0 myNMOS l=1u w=5u
V_DD N001 0 1.8
V_i+ N002 0 SINE(0.9 1m 1k)
V_i- N003 0 0.9
I1 N007 N004 20µ
