** sch_path: /home/nguyen2604/projects/DECODER3TO8/Schematic/CMOS_DECODER3_8.sch
**.subckt CMOS_DECODER3_8
x1 net4 Y0 net3 Y1 Y2 net1 Y3 GND Y4 Y5 Y6 Y7 net2 DECODER3_8
V1 net1 GND 1.8
V2 net2 GND PULSE(0 1.8 0 100p 100p 40n 80n)
V3 net3 GND PULSE(0 1.8 0 100p 100p 20n 40n)
V4 net4 GND PULSE(0 1.8 0 100p 100p 10n 20n)
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran 100p 100n
.save all
.control
    run
    plot v(E)
    plot v(Y0)
    plot v(Y1)
    plot v(Y2)
    plot v(Y3)
    plot v(Y4)
    plot v(Y5)
    plot v(Y6)
    plot v(Y7)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /home/nguyen2604/projects/DECODER3TO8/Schematic/DECODER3_8.sym # of pins=13
** sym_path: /home/nguyen2604/projects/DECODER3TO8/Schematic/DECODER3_8.sym
** sch_path: /home/nguyen2604/projects/DECODER3TO8/Schematic/DECODER3_8.sch
.subckt DECODER3_8 A0 Y0 A1 Y1 Y2 VDD Y3 VSS Y4 Y5 Y6 Y7 A2
*.ipin A0
*.ipin A1
*.ipin A2
*.iopin VDD
*.iopin VSS
*.opin Y0
*.opin Y1
*.opin Y2
*.opin Y3
*.opin Y4
*.opin Y5
*.opin Y6
*.opin Y7
x1 VDD A0 Y0 A1 Y1 Y2 Y3 VSS net1 DECODER2_4_E
x2 VDD A0 Y4 A1 Y5 Y6 Y7 VSS A2 DECODER2_4_E
x3 VDD A2 net1 VSS INVERTER
.ends


* expanding   symbol:  /home/nguyen2604/projects/DECODER3TO8/Schematic/DECODER2_4_E.sym # of pins=9
** sym_path: /home/nguyen2604/projects/DECODER3TO8/Schematic/DECODER2_4_E.sym
** sch_path: /home/nguyen2604/projects/DECODER3TO8/Schematic/DECODER2_4_E.sch
.subckt DECODER2_4_E VDD A0 Y0 A1 Y1 Y2 Y3 VSS E
*.ipin A0
*.ipin A1
*.ipin E
*.opin Y0
*.opin Y1
*.opin Y2
*.opin Y3
*.iopin VDD
*.iopin VSS
x1 VDD A0 net5 VSS INVERTER
x2 VDD A1 net6 VSS INVERTER
x3 VDD net5 net1 net6 VSS AND
x4 VDD A0 net2 net6 VSS AND
x5 VDD net5 net3 A1 VSS AND
x6 VDD A0 net4 A1 VSS AND
x7 VDD net1 Y0 E VSS AND
x8 VDD net2 Y1 E VSS AND
x9 VDD net3 Y2 E VSS AND
x10 VDD net4 Y3 E VSS AND
.ends


* expanding   symbol:  /home/nguyen2604/projects/DECODER3TO8/Schematic/INVERTER.sym # of pins=4
** sym_path: /home/nguyen2604/projects/DECODER3TO8/Schematic/INVERTER.sym
** sch_path: /home/nguyen2604/projects/DECODER3TO8/Schematic/INVERTER.sch
.subckt INVERTER VDD IN OUT VSS
*.ipin IN
*.opin OUT
*.iopin VDD
*.iopin VSS
XM2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
XM1 OUT IN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0 mult=1
+ m=1
.ends


* expanding   symbol:  /home/nguyen2604/projects/DECODER3TO8/Schematic/AND.sym # of pins=5
** sym_path: /home/nguyen2604/projects/DECODER3TO8/Schematic/AND.sym
** sch_path: /home/nguyen2604/projects/DECODER3TO8/Schematic/AND.sch
.subckt AND VDD A Y B GND
*.ipin A
*.ipin B
*.opin Y
*.iopin VDD
*.iopin GND
x1 VDD net1 A B GND NAND
x2 VDD net1 Y GND INVERTER
.ends


* expanding   symbol:  /home/nguyen2604/projects/DECODER3TO8/Schematic/NAND.sym # of pins=5
** sym_path: /home/nguyen2604/projects/DECODER3TO8/Schematic/NAND.sym
** sch_path: /home/nguyen2604/projects/DECODER3TO8/Schematic/NAND.sch
.subckt NAND VDD OUT IN1 IN2 VSS
*.ipin IN1
*.ipin IN2
*.opin OUT
*.iopin VDD
*.iopin VSS
XM1 OUT IN2 net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM2 net1 IN1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM3 OUT IN2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
XM4 OUT IN1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
.ends

.GLOBAL GND
.end
