magic
tech sky130A
timestamp 1762022518
<< nwell >>
rect 810 350 1045 515
<< nmos >>
rect 950 170 965 295
<< pmos >>
rect 950 370 965 495
<< ndiff >>
rect 890 275 950 295
rect 890 190 910 275
rect 930 190 950 275
rect 890 170 950 190
rect 965 275 1025 295
rect 965 190 985 275
rect 1005 190 1025 275
rect 965 170 1025 190
<< pdiff >>
rect 890 475 950 495
rect 890 390 910 475
rect 930 390 950 475
rect 890 370 950 390
rect 965 475 1025 495
rect 965 390 985 475
rect 1005 390 1025 475
rect 965 370 1025 390
<< ndiffc >>
rect 910 190 930 275
rect 985 190 1005 275
<< pdiffc >>
rect 910 390 930 475
rect 985 390 1005 475
<< psubdiff >>
rect 830 275 890 295
rect 830 190 850 275
rect 870 190 890 275
rect 830 170 890 190
<< nsubdiff >>
rect 830 475 890 495
rect 830 390 850 475
rect 870 390 890 475
rect 830 370 890 390
<< psubdiffcont >>
rect 850 190 870 275
<< nsubdiffcont >>
rect 850 390 870 475
<< poly >>
rect 950 495 965 510
rect 950 295 965 370
rect 950 155 965 170
rect 925 145 965 155
rect 925 125 935 145
rect 955 125 965 145
rect 925 115 965 125
<< polycont >>
rect 935 125 955 145
<< locali >>
rect 835 475 945 490
rect 835 390 850 475
rect 870 390 910 475
rect 930 390 945 475
rect 835 375 945 390
rect 970 475 1020 490
rect 970 390 985 475
rect 1005 390 1020 475
rect 970 375 1020 390
rect 995 290 1020 375
rect 835 275 945 290
rect 835 190 850 275
rect 870 190 910 275
rect 930 190 945 275
rect 835 175 945 190
rect 970 275 1020 290
rect 970 190 985 275
rect 1005 190 1020 275
rect 970 175 1020 190
rect 995 155 1020 175
rect 810 145 965 155
rect 810 130 935 145
rect 925 125 935 130
rect 955 125 965 145
rect 995 130 1045 155
rect 925 115 965 125
<< viali >>
rect 850 390 870 475
rect 910 390 930 475
rect 850 190 870 275
rect 910 190 930 275
<< metal1 >>
rect 810 475 1045 490
rect 810 390 850 475
rect 870 390 910 475
rect 930 390 1045 475
rect 810 375 1045 390
rect 810 275 1045 290
rect 810 190 850 275
rect 870 190 910 275
rect 930 190 1045 275
rect 810 175 1045 190
<< labels >>
rlabel locali 810 142 810 142 7 A
port 1 w
rlabel locali 1045 142 1045 142 3 Y
port 2 e
rlabel metal1 810 435 810 435 7 VP
port 3 w
rlabel metal1 810 235 810 235 7 VN
port 4 w
<< end >>
